module s1_control(
    
);

endmodule