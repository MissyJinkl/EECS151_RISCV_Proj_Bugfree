// TODO: change these paths if you move the Memory or RegFile instantiation
// to a different module
`define RF_PATH   cpu.rf
`define DMEM_PATH cpu.dmem
`define IMEM_PATH cpu.imem
`define BIOS_PATH cpu.bios_mem
`define CSR_PATH  cpu.tohost_csr
//`define CSR_PATH  cpu.csr_reg